LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY ALU IS
PORT(
  A, B : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  funct : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
  res : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END ALU;

ARCHITECTURE structural OF ALU IS

COMPONENT mux4to1 IS
PORT(
  a, b, c, d : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  s : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
  o1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

COMPONENT DIFF IS
PORT(
  i1, i2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  o1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

COMPONENT MULT IS
PORT(
  i1, i2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
  o1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

COMPONENT SUM IS
PORT(
  i1, i2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  o1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

COMPONENT CMP IS
PORT(
  i1, i2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  o1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

SIGNAL ssum, sdiff, smult, scmp : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
  unit0_0: SUM PORT MAP(A, B, ssum);
  unit0_1: DIFF PORT MAP(A, B, sdiff);
  unit0_2: MULT PORT MAP(A(3 DOWNTO 0), B(3 DOWNTO 0), smult);
  unit0_3: CMP PORT MAP(A, B, scmp);
  unit1: mux4to1 PORT MAP(ssum, sdiff, smult, scmp, funct, res);
END structural;
