LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY counter_tb IS
END counter_tb;

ARCHITECTURE arc OF counter_tb IS
COMPONENT counter IS
PORT(
  clock_enable, clock, reset: IN STD_LOGIC;
  outpt: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END COMPONENT;

SIGNAL clock_enable, clock, reset : STD_LOGIC;
SIGNAL outpt : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
  test_unit: counter PORT MAP(clock_enable, clock, reset, outpt);
  PROCESS
  BEGIN
    reset <= '1';
    WAIT FOR 10 ps;
    reset <= '0';
    WAIT FOR 10 ps;
    clock_enable <= '0';

    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;
    clock <= '1';
    WAIT FOR 10 ps;
    clock <= '0';
    WAIT FOR 10 ps;

  END PROCESS;
END arc;
